module uart_tb();
  
bit        PCLK_TB;
bit        PCLKG_TB;
bit        PRESETn_TB;
bit        PSEL_TB;
bit [11:2] PADDR_TB;
bit        PENABLE_TB;
bit        PWRITE_TB;
bit [31:0] PWDATA_TB;
bit [3:0]  ECOREVNUM_TB;
bit        RXD_TB;
bit [31:0] PRDATA_TB;
bit        PREADY_TB;
bit        PSLVERR_TB;
bit        TXD_TB;
bit        TXEN_TB;
bit        BAUDTICK_TB;
bit        TXINT_TB;
bit        RXINT_TB;
bit        TXOVRINT_TB;
bit        RXOVRINT_TB;
bit        UARTINT_TB;


 ////////////////////INSTANTIATION////////////////////

 cmsdk_apb_uart DUT (
 .PCLK(PCLK_TB),
 .PCLKG(PCLKG_TB),
 .PRESETn(PRESETn_TB),
 .PSEL(PSEL_TB),
 .PADDR(PADDR_TB),
 .PENABLE(PENABLE_TB),
 .PWRITE(PWRITE_TB),
 .PWDATA(PWDATA_TB),
 .ECOREVNUM(ECOREVNUM_TB),
 .PRDATA(PRDATA_TB),
 .PREADY(PREADY_TB),
 .PSLVERR(PSLVERR_TB),
 .RXD(RXD_TB),
 .TXD(TXD_TB),
 .TXEN(TXEN_TB),
 .BAUDTICK(BAUDTICK_TB),
 .TXINT(TXINT_TB),
 .RXINT(RXINT_TB),
 .TXOVRINT(TXOVRINT_TB),
 .RXOVRINT(RXOVRINT_TB),
 .UARTINT(UARTINT_TB)
 );


 
////////////////////CLOCK GENERATION////////////////////

localparam  CLK_PERIOD=10 ;

always #(CLK_PERIOD/2)  PCLK_TB = ~PCLK_TB ;
always #(CLK_PERIOD/2)  PCLKG_TB = ~PCLKG_TB ;

////////////////////INTERNAL REGISTER ADDRESS////////////////////

localparam [9:0] DATA = 10'h0;
localparam [9:0] STATE = 10'h1;
localparam [9:0] CTRL = 10'h2;
localparam [9:0] INTCLEAR = 10'h3;
localparam [9:0] INTSTATUS = 10'h3;
localparam [9:0] BAUDDIV = 10'h4;




////////////////////INITIALIZATION////////////////////

task initialize ;
begin
  PCLK_TB<= 0;
  PCLKG_TB<= 0;
  PSEL_TB<= 0; 
  PADDR_TB<= 0;
  PENABLE_TB<= 0;
  PWRITE_TB<= 0;
  ECOREVNUM_TB<= 0;
  PWDATA_TB<= 0;
  RXD_TB<= 1;
end
endtask


////////////////////RESET////////////////////

task reset;
begin
    PRESETn_TB <= 1'b0;
    #(CLK_PERIOD*10);
    PRESETn_TB <= 1'b1;
    #(CLK_PERIOD*10);
end
endtask

////////////////////TRANSFER USING APB TRANSFER////////////////////

task APB_TRANS ;
input [9:0] address;
input write ;
input [31:0] data;
begin
    @(posedge PCLK_TB)
    PADDR_TB <= address;
    PWRITE_TB <= write;
    PWDATA_TB <= data;
    PSEL_TB <= 1'b1;
    PENABLE_TB <= 1'b0;
    @(posedge PCLK_TB)
    PENABLE_TB <= 1'b1;
end
endtask

////////////////////RECEIVE////////////////////

task receive ;
  input [9:0] data ;
  int i;
  begin
    @(posedge PCLK_TB)
    PADDR_TB <= DATA;
    PSEL_TB <= 1;
    PENABLE_TB <=0;
    PWRITE_TB <= 0;
    for (i = 0 ; i < 10 ; i = i+1)
    begin
      RXD_TB = data[i] ;
      repeat(16)
      @(posedge PCLK_TB);
    end
    
  end
endtask





initial
begin
  
$dumpfile("uart.vcd") ;       
$dumpvars; 
initialize();
reset();
#(CLK_PERIOD*10);

APB_TRANS(CTRL,1,10'b111101);

APB_TRANS(DATA,1,8'b11010010);
APB_TRANS(DATA,1,8'b10010010);
repeat(7)
@(posedge PCLK_TB);
APB_TRANS(INTCLEAR,1,4'b0001);
repeat(7)
@(posedge PCLK_TB);
APB_TRANS(DATA,1,8'b10101001);
repeat(7)
@(posedge PCLK_TB);
APB_TRANS(INTCLEAR,1,1'b1);
APB_TRANS(DATA,1,8'b11101101);
repeat(50)
@(posedge PCLK_TB);

APB_TRANS(CTRL,1,10'b111110);

receive(10'b1100100100);

APB_TRANS(CTRL,1,10'b111111);
repeat(10)
@(posedge PCLK_TB);
fork
  begin
    APB_TRANS(DATA,1,10'b10010111);
  end
  begin
repeat(4)
@(posedge PCLK_TB);
    receive(10'b1010110100);
  end

join

#(1000*CLK_PERIOD);
$stop;
end

endmodule







